// module our_relay(o)